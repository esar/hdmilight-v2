
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package prog_mem_content is

-- content of p_0 ----------------------------------------------------------------------------------
constant p0_00 : BIT_VECTOR := X"C002E0E0E6A0BFCDE0D4BE1FC01BC01DC01FC021C023C025C027C029C02BC012";
constant p0_01 : BIT_VECTOR := X"0FE82FE201C0C007E0E081AA306393DFCFD1D1EE07B1921DE0B1E01107B1920D";
constant p0_02 : BIT_VECTOR := X"93DF950891DFE090C002E680E0F023229611539024110293E03A81BDF7B1912C";
constant p0_03 : BIT_VECTOR := X"B7CDE783B7FED000D000912CE0B02322963153A0241102A3E03A2DE080023062";
constant p0_04 : BIT_VECTOR := X"E04A2DE08002F00901FC91CFD20CE78ABF8DBF9EB60FB79ED513832483B3839A";
constant p0_05 : BIT_VECTOR := X"BF8DBF9EB60FB79EB548E08ABD87B568E0889530273323339631532024110224";
constant p0_06 : BIT_VECTOR := X"D1C0E982BF8DBF9EB60FB79ED4C78740835683648333938E9612B7ADE884B7FE";
constant p0_07 : BIT_VECTOR := X"C00924FF91FC961423229631531024110213E03A971391EDC0663064931F92FF";
constant p0_08 : BIT_VECTOR := X"D531D4DF23229631530024110203E03A971791EDF7A181200EF82EF924110243";
constant p0_09 : BIT_VECTOR := X"821582139711939CB7BEE0909631B7EDBE0F94F8970AB78DD529D52BD4D9D52F";
constant p0_0A : BIT_VECTOR := X"971391EDC0583064931F92FF90FF911FE090C003BE0F94F8960AB78D86118217";
constant p0_0B : BIT_VECTOR := X"F7B181200F082F0201C0C007E00091FC9614232296310EF2ED4001C02D4FE03A";
constant p0_0C : BIT_VECTOR := X"D0002F18E090D4B7D465D4BBD4BDD46B23229631531024110213E03A971791ED";
constant p0_0D : BIT_VECTOR := X"931F92FF92DF90FF911FE090C003900F900F82139711939CB7BEE0909631B7ED";
constant p0_0E : BIT_VECTOR := X"F35032C083005FEAF049300D0511D0B0F3D13F0F018CE0D0C002E0C02EE993DF";
constant p0_0F : BIT_VECTOR := X"01FC939C4F9E01C9238832804F3F921195702777E050E03001D92D9E82185FCA";
constant p0_10 : BIT_VECTOR := X"92DF92BF950890EF910F91CF2F844FFE01F9075796125F4F2388F01981805F2F";
constant p0_11 : BIT_VECTOR := X"2ED52EC51CF194082EB62EA6D396E090D06BE881BE0F94F89760B7CD93DF92FF";
constant p0_12 : BIT_VECTOR := X"C01134893583358281FAF754900FD34982D2B7ED2F18E068900FD35582B2B7ED";
constant p0_13 : BIT_VECTOR := X"2F61CFC22F61CFC6F641F021F0518181DDEE01C7DDC401C7DE2F01C7F6E1F039";
constant p0_14 : BIT_VECTOR := X"95089380939001C92F28C003EF2FFC009508E090CFFDB400DFFAF4112F18CFBE";
constant p0_15 : BIT_VECTOR := X"971191ED950891DF019CE08A238891F091E09509C00CEF2F2B899190918093DF";
constant p0_16 : BIT_VECTOR := X"9508932E96155F2F1FF3F44C1728919C9616913C9614973091FC96129509F019";
constant p0_17 : BIT_VECTOR := X"F04C070A16E881AE818C810A80E805710551F121859E01E993DF931F92FF92DF";
constant p0_18 : BIT_VECTOR := X"926F924F922F90CF90EF910F91CFF37C070A16E881AE818C1D011CE1DFB801C6";
constant p0_19 : BIT_VECTOR := X"920DE181EFE401DE0169012CBE0F94F897E1B7CD93DF930F92EF92CF92AF928F";
constant p0_1A : BIT_VECTOR := X"01B71E9D2C91E1922422017A2C31E0210B061AE424FFC00BF46904C116A8F7E1";
constant p0_1B : BIT_VECTOR := X"9381E28D2823051104F1018D01DAD36B019501C8938D81800FE60FECE0E101A6";
constant p0_1C : BIT_VECTOR := X"E070E050F4218990E070E05083B3839101F3E0A01B8E01CD200001DF01FE01D4";
constant p0_1D : BIT_VECTOR := X"94F896E101932F76FD57895001F3051F4010DF0E01D8C0040EEC2EE801840193";
constant p0_1E : BIT_VECTOR := X"92BF929F927F925F923F9508903F905F907F909F90BF90DF90FF911F91CFBE0F";
constant p0_1F : BIT_VECTOR := X"861F01C432651C5194082C31E0E1017ABFCDBFDEB60FB7DE93CF931F92FF92DF";
constant p0_20 : BIT_VECTOR := X"1461F0085380916C1CB194082E67C003246624CC87AB8789E0A0EF8FE2808A19";
constant p0_21 : BIT_VECTOR := X"1CB194081F4A0F2895A027AA9590279901ACD290E040E02A01CAE050E030F149";
constant p0_22 : BIT_VECTOR := X"9590279901ACD264E040E02A01CAE050E030876D3360875C873AF30853808110";
constant p0_23 : BIT_VECTOR := X"27335481CF9908A1862E8758833EF3085380911C1CB194081F4A0F2895A027AA";
constant p0_24 : BIT_VECTOR := X"C0BA0591C026F009F13132850591CF800591F4BC3685059101C99680F4189530";
constant p0_25 : BIT_VECTOR := X"E265CF572EC6C02FF0093788F4093783C0C80591F42C3781F4093780C0D40591";
constant p0_26 : BIT_VECTOR := X"2F76FD57915C01D70CCE2EC4C00C816281401CDF2CD1E054346428CD8A28C0B6";
constant p0_27 : BIT_VECTOR := X"F7E9900D911C01D7E030E01001C4816281401CDF2CD1E03401760172E020E00A";
constant p0_28 : BIT_VECTOR := X"01D801C49161C0050192E070E050F4218999E070E05083BC839AE0B00B919701";
constant p0_29 : BIT_VECTOR := X"1B8001CD200001D80EEEE0E205B197001DA187BC879A09B1970185AB85892388";
constant p0_2A : BIT_VECTOR := X"F491F41CF069C01EDD6401F74F1F0187DD9001C495602766894883AB8389E0A0";
constant p0_2B : BIT_VECTOR := X"CE7B236601D51CA1CE9D1CA1DD48C00101C4E06DC00701C4E067C0063762366E";
constant p0_2C : BIT_VECTOR := X"9728B7CD93DF902F904F906F908F90AF90CF90EF910F91DFBFCDBFDEB60FE090";
constant p0_2D : BIT_VECTOR := X"019C01A9856D01CE8618821E821C839A5F21C012E020970091909180BE0F94F8";
constant p0_2E : BIT_VECTOR := X"B5832F322F542B4A2B28E0A0B5842F322F54E040B525950891CFBE0F94F89628";
constant p0_2F : BIT_VECTOR := X"BD89B589BF81B781708C950801B92B4A2B28E0A0B5822F322F542B4A2B28E0A0";
constant p0_30 : BIT_VECTOR := X"9601E090BD89B58905919601E090BD89B589E081FC02F7D9308A0000E0807F87";
constant p0_31 : BIT_VECTOR := X"E0807F8BF7D9308A0000E0806088BD89B589E08005919601E090BD89B5890591";
constant p0_32 : BIT_VECTOR := X"0000000000006088C002B589FF372F38F7D9308A0000E0807F87F7D9308A0000";
constant p0_33 : BIT_VECTOR := X"0000E0807F8BBD89B5890F3330280000000000006084F7D9308A0000E0807F8B";
constant p0_34 : BIT_VECTOR := X"E090BD89B589E0307081952A9596E090F7D1302A5F2FE030BD89B589F7D9308A";
constant p0_35 : BIT_VECTOR := X"01D09508F6F95F3F05919601E090BD89B5897081954A9596E090B78005919601";
constant p0_36 : BIT_VECTOR := X"1BAAE2A1241101BD1DE19F631DE19F720DF00DF00DF00DF01DF19F640DE001F0";
constant p0_37 : BIT_VECTOR := X"94F801CF01AC95909570F7691F991F770BF50BB3F02007E417A21FEE1FAA01FD";
constant p0_38 : BIT_VECTOR := X"250067693A72000A20646425642564643A72000A3D6465757620646172724B4F";
constant p0_39 : BIT_VECTOR := X"316C2031646172720A643A645200617672642031762064643A72000A3D646425";
constant p0_3A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFF000044433938353431303E0A203E213841006464";
constant p0_3B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant p0_3C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant p0_3D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant p0_3E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant p0_3F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of p_1 ----------------------------------------------------------------------------------
constant p1_00 : BIT_VECTOR := X"9005E0FEE0B0E011BFDEE5CF2411C01CC01EC020C022C024C026C028C02AC02C";
constant p1_01 : BIT_VECTOR := X"961153E0241102E3E03A81BBF51901EC93CFC6D0F7E132A8C001E0A6F7D930A6";
constant p1_02 : BIT_VECTOR := X"01FC93CF91CFD245E683E090A390F7B1912C0F982F9201C0C007E09081AC2322";
constant p1_03 : BIT_VECTOR := X"B7DEE0909631B7EDD00097909690F7B181200FA82FA201C0C007E0A081F3F571";
constant p1_04 : BIT_VECTOR := X"C007E02081F3C0423062950891DFE090C003BE0F94F89606B78D821583A28389";
constant p1_05 : BIT_VECTOR := X"B7EDBE0F94F8970AB78DBD87B558E089BD87BD26FD27F7B181300F282F2301C0";
constant p1_06 : BIT_VECTOR := X"9508E0909508BE0F94F8960AB78D86118217821583229711939CB7BEE0909631";
constant p1_07 : BIT_VECTOR := X"2D4FE03A971591EDF7B181200F182F1201C0C007E01091FC9612F00901DC930F";
constant p1_08 : BIT_VECTOR := X"2D8F2F81F7B181200F082F0201C0C007E00091FC9616232296310EF2ED9001C0";
constant p1_09 : BIT_VECTOR := X"831682F48312938E9612B7ADE98DB7FEBF8DBF9EB60FB79ED5062F802F81D50C";
constant p1_0A : BIT_VECTOR := X"24FF91FC9612F00901DC930F9508910FD14FEA8ABF8DBF9EB60FB79ED4568700";
constant p1_0B : BIT_VECTOR := X"961623229631530024110203E03A971591EDF7A181200EF82EF424110243C009";
constant p1_0C : BIT_VECTOR := X"D000D490D4FCE0802F81D4982F802D8FF7B181200F182F1201C0C007E01091FC";
constant p1_0D : BIT_VECTOR := X"93CF930F92EF9508910FD0E9EC8F900F900FD3EC8312938E9612B7ADEC85B7FE";
constant p1_0E : BIT_VECTOR := X"CFE705D196214FFE01FE0511F061300A2F800718EF8FD0C5E1CFE0D02ED62EF8";
constant p1_0F : BIT_VECTOR := X"C002938E96115F8AF0D1F3D181805F2FC01BFD672D6DE040E020019C2D8F4FDE";
constant p1_10 : BIT_VECTOR := X"92EF92CF92AF90DF90FF911F91DFCFE15FEAF42417464F5FF7C1963132804F3F";
constant p1_11 : BIT_VECTOR := X"D000E050EE5F1CE1017EE060EE6BD06DEE85E092BFCDBFDEB60FB7DE93CF931F";
constant p1_12 : BIT_VECTOR := X"3587F709F41CF051818081E91611900F82C1B7FED000DF7001C7900F82A1B7FE";
constant p1_13 : BIT_VECTOR := X"DED401C7DE6401C7D37D348935873582CFCF2F61CFD32F61CFD72F61C0083588";
constant p1_14 : BIT_VECTOR := X"93CF012601279508E030B581EF3FC003B400911FE080FC03BD11E08D308A931F";
constant p1_15 : BIT_VECTOR := X"973091FC01DC91CF01C99509F7B90127012681889621EF3FF4290127012601EC";
constant p1_16 : BIT_VECTOR := X"92CF9714933C4F3F83600FE207399717918D9715912DF0A1971391ED95082F86";
constant p1_17 : BIT_VECTOR := X"C011071B06F981BF819D811B80F9F0F9056115412B89858D016C93CF930F92EF";
constant p1_18 : BIT_VECTOR := X"927F925F923F950890DF90FF911F91DF071B06F981BF819D1D111CF19408856C";
constant p1_19 : BIT_VECTOR := X"50819001E0F0961101370158BFCDBFDEB60FB7DE93CF931F92FF92DF92BF929F";
constant p1_1A : BIT_VECTOR := X"019501C80E8C2E892433018BC0042E220B170AF5018724EEFF7704D104B1E08A";
constant p1_1B : BIT_VECTOR := X"014F01F4F021F719050114E1017C01C901A601B7014D01D41FF71FFDE0F0D37A";
constant p1_1C : BIT_VECTOR := X"01C2E060E0412B898587E060E04083A28380E0B00B9F9701F7E9900D9672921C";
constant p1_1D : BIT_VECTOR := X"BFDEB60FDF2301C2956027668547F7B8150E5001916C01C21EFD2CF1E182DF3D";
constant p1_1E : BIT_VECTOR := X"92CF92AF928F926F924F922F902F904F906F908F90AF90CF90EF910F91DFBFCD";
constant p1_1F : BIT_VECTOR := X"861EC0C1F011C1801C41012E2E2E015B014CBE0F94F89761B7CD93DF930F92EF";
constant p1_20 : BIT_VECTOR := X"0471C05D308A2F8601D51CA12C71E071247724DD87BC879AE0B0E79F878D8A18";
constant p1_21 : BIT_VECTOR := X"01F51CA11F5B1F392FBAFD9797C0FD872F81019BE050E03001B9C019E040E020";
constant p1_22 : BIT_VECTOR := X"97C0FD872F81019BE050E03001B9C019E040E020F409C02D874B8729308A2F81";
constant p1_23 : BIT_VECTOR := X"FD272F262F8608B19408863F834F832D308A2F8101D51CA11F5B1F392FBAFD97";
constant p1_24 : BIT_VECTOR := X"3683F409358CC0DD978D0591F43C328FF409328E0591F1D13684C00101C9318A";
constant p1_25 : BIT_VECTOR := X"DDFB01C42CD1E061C0BF0591C0440591C009F009368C0591C0400591C0ACF009";
constant p1_26 : BIT_VECTOR := X"01C495602766914D1CDF2CD1E0428173815101F70CCE2EC5F459F411CF508A39";
constant p1_27 : BIT_VECTOR := X"01CD200001D8910DCFECE020E1008173815101F70CCE2EC3C08FDE34E030E010";
constant p1_28 : BIT_VECTOR := X"918CDD9D018F01F8DDC701C4E060E0412B898988E060E04083AB8389E0A01B80";
constant p1_29 : BIT_VECTOR := X"0B919701F7E9900D1EFFE0F0F72905A11DB1960187AB878909A185BC859AF091";
constant p1_2A : BIT_VECTOR := X"C0053661366936680178816001C45F0CC02701922F76FD57895983BC839AE0B0";
constant p1_2B : BIT_VECTOR := X"E080F009916C1CB194081CB1940801C4E06AC00401C4E068C00A01C4F469F061";
constant p1_2C : BIT_VECTOR := X"B60FB7DE93CF9508903F905F907F909F90BF90DF90FF911F91CFBE0F94F89661";
constant p1_2D : BIT_VECTOR := X"01C9DE17857E9601821F821D821B83894F3F019EE030F41901270126BFCDBFDE";
constant p1_2E : BIT_VECTOR := X"E09027222F432B5B2B39E0B0E09027222F43E050E030BC1291DFBFCDBFDEB60F";
constant p1_2F : BIT_VECTOR := X"B5897F8B9508708CBD89B58901CA2B5B2B39E0B0E09027222F432B5B2B39E0B0";
constant p1_30 : BIT_VECTOR := X"308A0000E0806084F7D9308A0000E08060889508C002B60005919601E090BD89";
constant p1_31 : BIT_VECTOR := X"E090BD89B58905919601E090BD89B58960849508F7D9308A0000E0807F87F7D9";
constant p1_32 : BIT_VECTOR := X"B58900000000BD89B5897F87C003E020950805919601E090BD89B58905919601";
constant p1_33 : BIT_VECTOR := X"9601E090BD89B5897F87CFDCF0115F2F00000000BD89B58905919601E090BD89";
constant p1_34 : BIT_VECTOR := X"0000E0807F8BE0209508F7E19587E0232F8905314F3F0000E0206084B7900591";
constant p1_35 : BIT_VECTOR := X"9F739F622F823038F7D9308A0000E08060842B28F7E19587E0430F22F7D9308A";
constant p1_36 : BIT_VECTOR := X"1BBB2E1A950801CF1FF90DB01FF90DB027999F659F749F839F920DE01DF19F82";
constant p1_37 : BIT_VECTOR := X"CFFF950801BD019B95809560941A1F881F660BE41BA207F507B31FFF1FBBC00D";
constant p1_38 : BIT_VECTOR := X"3D6474686C20726564252520203A007261207265642525006C617264203A6500";
constant p1_39 : BIT_VECTOR := X"612061767264203A650025206165326C203264616C6131726120726564252520";
constant p1_3A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF464542413736333200200D000A0052563272";
constant p1_3B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant p1_3C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant p1_3D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant p1_3E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant p1_3F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

end prog_mem_content;

